(************************************)
(*                                  *)

         module "Mld_hash"

(*                                  *)
(************************************)

" <hash> : Set hash type you want to compute (ed2k, sig2dat,bp)" = " <hash> : Set hash type you want to compute (ed2k, sig2dat,bp)"

" <nth size>: check C file functions" = " <nth size>: check C file functions"

" <filenames> : compute hashes of filenames" = " <filenames> : compute hashes of filenames"

(************************************)
(*                                  *)

         module "Former Translation"

(*                                  *)
(************************************)

"Misc" = "\214vrigt"

"Client" = "Klient"

"GUI" = "Anv\228ndargr\228nssnitt"

"Columns titles" = "Kolumntitlar"

"Shared files upload info" = "Uppladdningsinfo f\246r delade filer"

"Columns for the results of searches and files of a friends" = "Kolumner f\246r resultat efter s\246kningar efter s\246kningar efter filer"

"Columns for the locations of a file" = "Kolumner f\246r filplatser"

"File locations" = "Filplatser"

"Columns for the friends" = "Kolumner f\246r v\228nner"

"Columns for the downloaded files" = "Kolumner f\246r nedladdade filer"

"Columns for the files being downloaded" = "Kolumner f\246r filer under nedladdning"

"Columns for the servers" = "Kolumner f\246r servrar"

"Style of toolbars" = "Typ av verktygsf\228lt"

"What is displayed in toolbar buttons : text, icon or both" = "Hur visas verktygsf\228ltets knappar: text, ikon eller b\229da?"

"Use relative %% availability" = "Anv\228nd relativ %% tillg\228nglighet"

"Calculate %% availability ignoring already present chunks" = "Ber\228kna %% tillg\228nglighet utan nedladdade stycken"

"Display the availability of a chunk as height or color coded bar" = "Visa tillg\228ngigheten f\246r stycken som h\246jd eller f\228rgkodad stapel"

"Use size suffixes (G, M, k)" = "Anv\228nd storlekssuffix (G, M, k)"

"Auto-resize lists columns" = "Automatisk storkleksinst\228llnig f\246r kolumner"

"Auto-resize" = "Automatisk storkleksinst\228llnig"

"Colors" = "F\228rger"

"Files listed" = "Listade filer"

"Color for not connected servers or users" = "F\228rg f\246r ej anslutna servrar och anv\228ndare"

"Color for connected servers or users" = "F\228rg f\246r anslutna servrar och anv\228ndare"

"Color for unavailable files" = "F\228rg f\246r filer som ej \228r tillg\228ngliga"

"Not available" = "Ej tillg\228ngliga"

"Color for available files, not downloading" = "F\228rg f\246r tillg\228ngliga filer som inte laddas ner"

"Available" = "Tillg\228nglig"

"Color for files being downloaded" = "F\228rf f\246r filer som laddas ner"

"Color for downloaded files" = "F\228rg f\246r nedladdade filer"

"Default color in lists" = "Standardf\228rg i listor"

"Default" = "Standard"

"GUI server" = "Anv\228ndargr\228nssnittsserver"

"The password to use when connecting to the server" = "L\246senord att anv\228nda vid anslutning till server"

"The server hostname to connect to" = "Serverv\228rdnamn att ansluta till"

"Hostname" = "V\228rdnamn"

"The server port to connect to" = "Serverport att ansluta till"

"Extended Search" = "Ut\246kad s\246kning"

"Local Search" = "S\246k lokalt"

"Comment" = "Kommentar"

"Track number" = "L\229tnummer"

"Year" = "\197r"

"Rooms" = "Rum"

"Results" = "Resultat"

"Queries" = "Fr\229gor"

"Settings" = "Inst\228llningar"

"Help" = "Hj\228lp"

"Quit" = "Avsluta"

"Reconnect" = "\197teranslut"

"Kill core" = "Avsluta k\228rna"

"File" = "Fil"

"Refresh" = "Uppdatera"

"Uploaded" = "Uppladdat"

"Uploads stats" = "Uppladdningsstatistik"

"Requests" = "F\246rfr\229gningar"

"Uploads" = "Uppladdningar"

"Show hidden fields" = "Visa dolda f\228lt"

"Browse files" = "Bl\228ddra filer"

"Display all servers" = "Visa alla"

"Remove all friends" = "T\246m"

"Find friend" = "Hitta v\228n"

"Get format info" = "Formatinfo"

"Preview" = "F\246rhandsvisa"

"Verify chunks" = "Verifiera delar"

"Pause/Resume" = "Pausa/Forts\228tt"

"Upload" = "Uppladdning"

"Direct" = "Direkt"

"Edit mp3 tags" = "Editera mp3-tags"

"Save file as" = "Spara fil som"

"Unknown" = "Ok\228nd"

"Done" = "Klar"

"Paused" = "Pausad"

"Cancelled" = "Avbruten"

"Downloading" = "Laddar ner"

"Queued" = "I k\246"

"Removed" = "Borttagen"

"Connected" = "Ansluten"

"Initiating" = "Initierar"

"Connecting" = "Ansluter"

"No" = "Nej"

"Yes" = "Ja"

"Kind" = "Slag"

"Clear Console" = "T\246m konsol"

"Console" = "Konsol"

"Command" = "Kommando"

"Set Option" = "St\228ll in"

"Value:" = "V\228rde:"

"Option:" = "Inst\228llning:"

"Client hostname" = "Klientens v\228rdnamn"

"Features" = "Finesser"

"Max Hits" = "Max tr\228ffar"

"Max server age (days)" = "Max server\229lder (dagar)"

"Remove old\nservers" = "Gallra"

"Recover MD4:" = "\197tervinn MD4:"

"Save" = "Spara"

"Save all" = "Spara allt"

"%d Downloaded Files" = "%d nedladdade filer"

"Downloaded Files: %d/%d" = "Nedladdade filer: %d/%d"

"Downloading Files" = "Filer att ladda ner"

"Connect" = "Anslut"

"Users" = "Anv\228ndare"

"Connect more\nservers" = "Fler servrar"

"Add friend" = "L\228gg till v\228n"

"Add server" = "L\228gg till server"

"Add to friends" = "L\228gg till bland v\228nner"

"Connected to %d / %d locations" = "Ansluten till %d / %d platser"

"Disconnect all" = "Koppla fr\229n alla"

"Retry connect" = "\197teranslut"

"Availability" = "Tillg\228nglighet"

"Downloaded" = "Nedladdade"

"Subscribe" = "Prenumerera"

"Force Download" = "Tvinga nedladdning"

"Download" = "Ladda ner"

"Download selected directory" = "Ladda ner vald mapp"

"Download selected files" = "Ladda ner valda filer"

"Properties" = "Egenskaper"

"Size" = "Storlek"

"Filename" = "Filnamn"

"Files" = "Filer"

"View users" = "Kolla v\228nner"

"View files" = "Kolla filer"

"Close room" = "L\228mna room"

"Remove" = "Ta bort"

"%d Results" = "%d Resultat"

"Submit" = "Skicka"

"Mp3 options" = "Mp3-inst\228llningar"

"Close" = "St\228ng"

"Stop" = "Avbryt s\246kning"

"Min bitrate" = "Minsta bitrate"

"Title" = "Titel"

"Browse" = "Bl\228ddra"

"Friend" = "V\228n"

"Type" = "Typ"

"Network" = "N\228tverk"

"Max size" = "St\246rsta storlek"

"Min size" = "Minsta storlek"

"Search" = "S\246kning"

"Query" = "Fr\229ga"

"Apply and save options" = "Aktivera och spara inst\228llningar"

"Client connection" = "Clientanslutning"

"Server connection" = "Serveranslutning"

"Upload limit (kB/s)" = "Uppladdningsbegr\228nsning (kB/s)"

"Download limit (kB/s)" = "Nedladdningsbegr\228nsning (kB/s)"

"Disconnect" = "Koppla fr\229n"

"Max connected clients" = "Max anslutna klienter"

"Max connected servers" = "Max anslutna servrar"

"Name" = "Namn"

"General" = "Generell"

"Gui refresh delay" = "Anv\228ndargr\228nssnittets uppdateringsf\246rdr\246jning"

"Long retry delay" = "L\229ng \229terf\246rs\246ksf\246rdr\246jning"

"Medium retry delay" = "Mellanstor \229terf\246rs\246ksf\246rdr\246jning"

"Small retry delay" = "Liten \229terf\246rs\246ksf\246rdr\246jning"

"Check serverDB connection" = "Kolla serverDB-anslutning"

"Check server connection" = "Kolla server-anslutning"

"Check client connections" = "Kolla klient-anslutningar"

"Save options delay" = "F\246rdr\246jning spara inst\228llningar"

"Delays" = "F\246rdr\246jningar"

"Ports" = "Portar"

"GUI port" = "Anv\228ndargr\228nssnittsport"

"Control port" = "Kontrollport"

"Connection port" = "Anslutningsport"

"No current search" = "Ingen p\229g\229ende s\246kning"

"Downloading %d file(s)" = "Laddar ner %d file(r)"

"Connected to %d/%d server(s)" = "Ansluten till %d/%d server/sevrar"

"Not connected" = "Ej ansluten"

"Options" = "Inst\228llningar"

"Searches" = "S\246kningar"

"Friends" = "V\228nner"

"Downloads" = "Nedladdnigar"

"Servers" = "Servrar"

"State" = "Tillst\229nd"

"Last seen" = "Senast sedd"

"Age" = "\197lder"

"Rate" = "Hastighet"

"Address" = "Adress"

"Password" = "L\246senord"

"Cancel" = "Avbryt"

