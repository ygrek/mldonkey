(*
 translated by kokamomi@gueststars.net
 s� det s�.
 
 Installation:
 # cp ~/.mldonkey_gui_messages.ini .mldonkey_gui_messages.ini.bak
 # cp /s�kv�g/till/din/mldonkey-distribution/i18n/gui_messages.ini.sv ~/.mldonkey_gui_messages.ini
 
*)

 ok = Ok
 cancel = Avbryt
 password = L�senord
 address = Adress
 percent = "%%"
 rate = Hastighet
 age = �lder
 last_seen = "Senast sedd"
 eta = "Tid kvar"
 priority = Prioritet
 state = Tillst�nd
 servers = Servrar
 downloads = Nedladdningar
 friends = V�nner
 searches = S�kningar
 options = Inst�llningar
 not_connected = "Ej ansluten"
 black_listed = "Svartlistade"
 connected_to_servers = "Ansluten till %d/%d server/sevrar"
 downloading_files = "Laddar ner %d file(r)"
 no_current_search = "Ingen p�g�ende s�kning"
 connection_port = "Anslutningsport"
 control_port = "Kontrollport"
 gui_port = "Anv�ndargr�nssnittsport"
 ports = Portar
 delays = F�rdr�jningar
 save_options_delay = "F�rdr�jning spara inst�llningar"
 check_client_connections = "Kolla klient-anslutningar"
 check_server_connection = "Kolla server-anslutning"
 check_serverDB_connection = "Kolla serverDB-anslutning"
 small_retry_delay = "Liten �terf�rs�ksf�rdr�jning"
 medium_retry_delay = "Mellanstor �terf�rs�ksf�rdr�jning"
 long_retry_delay = "L�ng �terf�rs�ksf�rdr�jning"
 gui_refresh_delay = "Anv�ndargr�nssnittets uppdateringsf�rdr�jning"
 general = Generell
 name = Namn
 max_connected_servers = "Max anslutna servrar"
 max_connected_clients = "Max anslutna klienter"
 disconnect = "Koppla fr�n"
 download_limit = "Nedladdningsbegr�nsning (kB/s)"
 upload_limit = "Uppladdningsbegr�nsning (kB/s)"
 timeouts = Timeouts
 server_connection = "Serveranslutning"
 client_connection = "Clientanslutning"
 save_and_apply_options = "Aktivera och spara inst�llningar"
 query = Fr�ga
 search = S�kning
 min_size = "Minsta storlek"
 max_size = "St�rsta storlek"
 media = Media
 format = Format
 network = N�tverk
 client_type = Typ
 album = Album
 friend = V�n
 contact = Bl�ddra
 artist = Artist
 title = Titel
 min_bitrate = "Minsta bitrate"
 stop_search = "Avbryt s�kning"
 close_search = "Avsluta s�kning"
 mp3_options = "Mp3-inst�llningar"
 submit = Skicka
 results = "%d Resultat"
 friends = V�nner
 ip = IP
 port = Port
 remove = "Ta bort"
 close = St�ng
 close_room = "L�mna room"
 view_files = "Kolla filer"
 view_users = "Kolla v�nner"
 files = Filer
 network = N�tverk
 display = Display
 filename = Filnamn
 size = Storlek
 properties = Egenskaper
 md4 = MD4
 download_selected_files = "Ladda ner valda filer"
 download_selected_dir = "Ladda ner vald mapp"
 download = "Ladda ner"
 force_download = "Tvinga nedladdning"
 subscribe = Prenumerera
 downloaded = Nedladdad
 availability = Tillg�nglighet
 cancel = Avbryt
 retry_connect = �teranslut
 disconnect_all = "Koppla fr�n alla"
 connected_to_locations = "Ansluten till %d / %d platser"
 add_to_friends = "L�gg till bland v�nner"
 add_server = "L�gg till server"
 add_friend = "L�gg till v�n"
 connect_more_servers = "Fler servrar"
 connect_more_servers_tips = "Anslut till fler servrar"
 users = Anv�ndare
 status = Status
 connect = Anslut
 disconnect = "Koppla fr�n"
 files_to_download = "Filer att ladda ner"
 downloaded_files = "Nedladdade filer: %d/%d"
 files_downloaded = "%d nedladdade filer"
 save_all = "Spara allt"
 save = Spara
 server_name = Name
 server_desc = Description
 server_nusers = Users
 server_nfiles = Files
 ed2k = "ed2k:"
 recover_md4 = "�tervinn MD4:"
 remove_old_servers = Gallra
 remove_old_servers_tips = "Gallra ut gamla servrar"
 max_server_age = "Max server�lder (dagar)"
 max_hits = "Max tr�ffar"
 features = Finesser
 hostname = "Klientens v�rdnamn"
 option_name = "Inst�llning:"
 option_value = "V�rde:"
 set_option = "St�ll in"
 command = Kommando
 console = Konsol
 clear_console = "T�m konsol"
 friend_kind = Slag
 friend_status = Status
 friend_name = Namn
 dialog = Chat
 yes = Ja
 no = Nej
 connecting = Ansluter
 initiating = Initierar
 connected = Ansluten
 removed = Borttagen
 queued = "I k�"
 downloading = "Laddar ner"
 cancelled = Avbruten
 paused = Pausad
 dl_done = Klar
 unknown = Ok�nd
 nusers = Anv�ndare
 save_as = "Spara fil som"
 edit_mp3 = "Editera mp3-tags"
 kind = Slag
 direct = Direkt
 upload = Uppladdning
 pause_resume_dl = "Pausa/Forts�tt"
 verify_chunks = "Verifiera delar"
 preview = F�rhandsvisa
 get_format = "Formatinfo"
 find_friend = "Hitta v�n"
 remove_all_friends = T�m
 remove_all_friends_tips = "Ta bort alla v�nner"
 toggle_display_all_servers = "Visa alla"
 toggle_display_all_servers_tips = "Visa alla servrar (�ven ej anslutna)"
 browse_files = "Bl�ddra filer"
 show_hidden_fields = "Visa dolda f�lt"
 uploads = Uppladdningar
 requests = F�rfr�gningar
 upstats = Uppladdningsstatistik
 uploaded = Uppladdat
 refresh = Uppdatera
 mFile = Fil
 mKill_server = "Avsluta k�rna"
 mFile = Fil
 mReconnect = �teranslut
 mDisconnect = "Koppla fr�n"
 mQuit = Avsluta
 mHelp = Hj�lp
 mSettings = Inst�llningar
 mServers = Servrar
 mDownloads = Nedladdningar
 mFriends = V�nner
 mConsole = Konsol
 mQueries = Fr�gor
 mResults = Resultat
 mRooms = Rum
 mUploads = Uppladdningar
 title = Titel
 artist = Artist
 album = Album
 year = �r
 tracknum = "L�tnummer"
 comment = Kommentar
 genre = Genre
 local_search = "S�k lokalt"
 extended_search = "Ut�kad s�kning"
 o_gui_port = "Anv�ndargr�nssnittsport"
 h_gui_port = "Serverport att ansluta till"
 o_hostname = V�rdnamn
 h_hostname = "Serverv�rdnamn att ansluta till"
 o_password = L�senord
 h_gui_password = "L�senord att anv�nda vid anslutning till server"
 o_gui_server = Anv�ndargr�nssnittsserver
 o_col_default = Standard
 h_col_default = "Standardf�rg i listor"
 o_col_downloaded = Nedladdade
 h_col_downloaded = "F�rg f�r nedladdade filer"
 o_col_downloading = "Laddar ner"
 h_col_downloading = "F�rf f�r filer som laddas ner"
 o_col_avail = Tillg�nglig
 h_col_avail = "F�rg f�r tillg�ngliga filer som inte laddas ner"
 o_col_not_avail = "Ej tillg�ngliga"
 h_col_not_avail = "F�rg f�r filer som ej �r tillg�ngliga"
 o_col_connected = Ansluten
 h_col_connected = "F�rg f�r anslutna servrar och anv�ndare"
 o_col_not_connected = "Ej ansluten"
 h_col_not_connected = "F�rg f�r ej anslutna servrar och anv�ndare"
 o_col_connecting = Ansluter
 o_col_files_listed = "Listade filer"
 o_colors = F�rger
 o_auto_resize = "Automatisk storkleksinst�llnig"
 h_auto_resize = "Automatisk storkleksinst�llnig f�r kolumner"
 o_files_auto_expand_depth = "Files auto-expand depth"
 o_use_size_suffixes = "Anv�nd storlekssuffix (G, M, k)"
 h_use_availability_height = "Visa tillg�ngigheten f�r stycken som h�jd eller f�rgkodad stapel"
 o_use_availability_height = "Use height encoded availability"
 h_use_relative_availability = "Ber�kna %% tillg�nglighet utan nedladdade stycken"
 o_use_relative_availability = "Anv�nd relativ %% tillg�nglighet"
 h_chunk_width = "Bredd p� segment i tilg�nlighetsstapeln"
 o_chunk_width = "Segmentbredd"
 h_toolbars_style = "Hur visas verktygsf�ltets knappar: text, ikon eller b�da?"
 o_toolbars_style = "Typ av verktygsf�lt"
 o_layout = Layout
 o_servers_columns = Servrar
 h_servers_columns = "Kolumner f�r servrar"
 o_downloads_columns = Nedladdnigar
 h_downloads_columns = "Kolumner f�r filer under nedladdning"
 o_downloaded_columns = Nedladdade
 h_downloaded_columns = "Kolumner f�r nedladdade filer"
 o_friends_columns = V�nner
 h_friends_columns = "Kolumner f�r v�nner"
 o_file_locations_columns = "Filplatser"
 h_file_locations_columns = "Kolumner f�r filplatser"
 o_results_columns = Resultat
 h_results_columns = "Kolumner f�r resultat efter s�kningar efter s�kningar efter filer"
 o_shared_files_up_colums = "Uppladdningsinfo f�r delade filer"
 o_columns = "Kolumntitlar"
 o_gui = Anv�ndargr�nssnitt
 o_client = Klient
 o_options = Inst�llningar
 o_misc = �vrigt

(*
 The following options are not used (errors, obsolete, ...) 
*)
